`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/13/2025 04:29:10 PM
// Design Name: 
// Module Name: fir_filter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module fir_filter(
input_data,clk,reset,enable,output_data,samplet
    );
    input clk,reset,enable;
    parameter n1=8,n2=16,n3=32;
    parameter numcoff=8;
    input signed [n2-1:0] input_data;
    output signed [n2-1:0] samplet;
    output signed [n3-1:0] output_data;
    wire signed [n1-1:0] b[0:7];

assign b[0] = 8'd16;
assign b[1] = 8'd16;
assign b[2] = 8'd16;
assign b[3] = 8'd16;
assign b[4] = 8'd16;
assign b[5] = 8'd16;
assign b[6] = 8'd16;
assign b[7] = 8'd16;

    
    reg signed [n3-1:0] output_data_reg;
    reg signed [n2-1:0] samples[0:6];
    
//    genvar i;
//    for(i=0;i<numcoff;i=i+1)
//    begin:bsvalue_assign
//    assign b[i]=8'b00010000;
//    end



    integer j;
    always @(posedge clk)
    begin
    if (reset)
    begin
    for(j=0;j<7;j=j+1)begin
    samples[j]<=0;end
     output_data_reg<=0;
    end
    if(enable &&(!reset)) begin
    output_data_reg<=b[0]*input_data+b[1]*samples[0]+b[2]*samples[1]+b[3]*samples[2]+b[4]*samples[3]
    +b[5]*samples[4]+b[6]*samples[5]+b[7]*samples[6];
    samples[0]<=input_data;
    for(j=1;j<7;j=j+1)begin
    samples[j]<=samples[j-1];
    end
    
    end
   
    end
    assign output_data=output_data_reg;
    assign samplet=samples[0];
endmodule
